netcdf {
  // Example 5
  // An aggregated data variable and an aggregated coordinate variable in the
  // same dataset. There are two external netCDF files, each of which contains a
  // fragment for each aggregation variable. The aggregation definition variables
  // for each aggregation variable are stored in different groups
  // (aggregation_temp and aggregation_time), but the file terms of the
  // aggregated_data attributes refer to a variable in the root group that stores
  // the external file names that apply to both aggregation variables.

  dimensions:
    // Aggregated dimensions
    time = 12 ;
    level = 1 ;
    latitude = 73 ;
    longitude = 144 ;
    // Fragment dimensions
    f_time = 2 ;
    f_level = 1 ;
    f_latitude = 1 ;
    f_longitude = 1 ;
    // Extra dimensions
    i = 4 ;
    ii = 1 ;
    j = 2 ;
  variables:
    // Data variable
    double temp ;
      temp:standard_name = "air_temperature" ;
      temp:units = "K" ;
      temp:cell_methods = "time: mean" ;
      temp:aggregated_dimensions = "time level latitude longitude" ;
      temp:aggregated_data = "location: /aggregation_temp/location
                              file: /aggregation_temp/aggregation_file
                              format: aggregation_format
                              address: /aggregation_temp/address" ;
    // Coordinate variables
    double time ;
      time:standard_name = "time" ;
      time:units = "days since 2001-01-01" ;
      temp:aggregated_dimensions = "time" ;
      temp:aggregated_data = "location: /aggregation_time/location
                              file: /aggregation_time/file
                              format: agregation_format
                              address: /aggregation_time/address" ;
    double level(level) ;
      level:standard_name = "height_above_mean_sea_level" ;
      level:units = "m" ;
    double latitude(latitude) ;
      latitude:standard_name = "latitude" ;
      latitude:units = "degrees_north" ;
    double longitude(longitude) ;
      longitude:standard_name = "longitude" ;
      longitude:units = "degrees_east" ;
    // Aggregation definition variables
    string aggregation_format ;

  // global attributes:
    :Conventions = "CF-1.9 CFA-0.6" ;
  data:
    temp = _ ;
    time = _ ;
    aggregation_format = "nc" ;

  group: aggregation_temp {
    variables:
      // Temperature aggregation definition variables
      int location(i, j) ;
      string file(f_time, f_level, f_latitude, f_longitude) ;
      string address(f_time, f_level, f_latitude, f_longitude) ;

    data:
      location = 6, 6,
                 1, _,
                 73, _,
                 144, _ ;
      file = "January-June.nc", "July-December.nc" ;
      address = "temp", "temp" ;
  }

  group: aggregation_time {
    variables:
      // Time aggregation definition variables
      int location(ii, j) ;
      string aggregation_file(f_time) ;
      string address(f_time) ;

    data:
      location = 6, 6 ;
      aggregation_file = "January-June.nc", "July-December.nc" ;
      address = "time", "time" ;
  }
}
